class my_test;

   top_final top_final();   

endclass // my_test
