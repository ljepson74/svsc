module asdf();

   initial begin
      repeat (33) $display("HI HO SILVER,  AWAY!");
   end
   
endmodule