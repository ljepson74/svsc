import uvm_pkg::*;

class env extends uvm_env;

   

endclass : env