lkj@srgo2img02.ba.imgtec.org.1196:1426158600