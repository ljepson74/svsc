module top;
   import uvm_pkg::*;
`include "uvm_macros.svh"

   initial begin
      run_test();
   end

endmodule : top
