class class_y;

   rand int int1;
   rand int int2;
   
/*   function new(input int one, two);
      int1=one;
      int2=two;
      $display(" new class_y and int1=%0d  int2=%0d",int1,int2);
   endfunction
  */ 

   function void show();
      $display("int1=%0d  int2=%0d",int1,int2);
   endfunction
endclass