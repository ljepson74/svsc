class class_stimulus;

   virtual 

   
endclass : class_stimulus
