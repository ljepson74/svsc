interface switch_interface(input clk);

   //your code here


endinterface
