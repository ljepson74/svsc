lkj@srgo2img02.ba.imgtec.org.22281:1441973250