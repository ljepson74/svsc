`include "packet.sv"

program testcase(...);

   //your code here
endprogram
