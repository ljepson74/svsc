//import branch_pkg::branch_hi;
import branch_pkg::*;

class trunk;
   function new();
      branch_hi();
      //leaf_hi();
   endfunction : new

endclass : trunk