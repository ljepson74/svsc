// TITLE: JOE IS LATE

// SECTION: LIANG IS GREAT
//  SECTION:  test1 extrawhitespace
// sECTION: test2 camcelcase LIANG IS GREAT
// section: test3 lowercase LIANG IS GREAT

// CLASS: TOP
class top();

   top2 m_top2;
endclass

