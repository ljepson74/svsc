class c2;
      
   function new(); 
      $display(" %m: MADE C2");      
   endfunction // new

   function void do_smthg;
      $display("RAAAR!  how was that?");      
   endfunction
   
endclass // c1
