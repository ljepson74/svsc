bind dut bound bound_u(.clk(clk), .data_bus(data_bus), .bus_data(bus_data));
