module cast;


endmodule : cast
