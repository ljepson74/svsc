interface my_if();
   logic  [7:0] some_data;
endinterface


     