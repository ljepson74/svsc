import uvm_pkg::*;

//class my_transaction extends uvm_sequence_item;
class a_transaction extends uvm_sequence;


/*
 function new(string name = "");
 super.new(name);
   endfunction: new
 */

endclass: a_transaction

