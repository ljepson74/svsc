module testbench();

   //your code here
endmodule
