module stimulus(
		score_items_if stimulus_if;
		);
   
   
   
endmodule // stimulus
