import uvm_pkg::*;
`include "uvm_macros.svh"

class svs_test extends uvm_test;
   `uvm_component_utils(svs_test)   
endclass : svs_test



   