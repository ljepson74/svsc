bind coin_counter assertion t2(clk,load,count,dispense,empty);

