interface score_if;

   integer if_age;
   integer if_iq;
   integer if_shoesize;
    
endinterface // score_if
