module irun_option_play;

   initial begin
      $display($time," Hey senoro");
      #113;      
      $display($time," Hey senoro");
      #5;      
      $display($time," Hey senoro");
      #7;      
      $display($time," Hey senoro");
      #9;      
   end
   

endmodule // irun_option_play
