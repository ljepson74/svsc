module top;


  initial begin
    $display(" this is a pretty long comment, but I will try to break it up \
a litlte bit more . %0s %0d","fredship",777, 
	     "how do you like that %0d %0d  %0d",1234, 5678, 91011121313);
    
  end
  
endmodule // top
