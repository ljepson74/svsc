lkj@srgo2img01.ba.imgtec.org.9303:1344457658