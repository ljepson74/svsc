package my_package1;

   import my_package2::*;
   
   int valueA;

   function void tellmex();
      $display("\n\n ***** bonjour ****\n\n");
   endfunction

endpackage : my_package1
