module top;

   initial begin
      $display("%m:  We are here");      
   end   

endmodule