module stimulus(
    output integer out_age,
    output integer out_iq,
    output integer out_shoesize
    );
    
    integer cnt;
/*    
    for (cnt=0; cnt<10; cnt++) begin
        #40ns;
        out_age = $urandom;
        out_iq  = $urandom;
        out_shoesize = $urandom;
    end 
  */  
    
endmodule   
    

