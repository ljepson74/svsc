interface d_if(
	       input logic clk
	       );

   logic [3:0] interface_bus;

endinterface