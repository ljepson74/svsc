/*
 Loose ideas for interview questions.
 
 a) Get the person in front of a terminal where they can work with real code.   It is too easy to hand-wave with pseudo-code
 
 */


////////////////////
////////////////////
//*) Array of objects.  Where objects are of simple class
//Does person know not just to new the array
array = new[5];
foreach (array[ii]) begin
   array[ii]=new();    //but to new each class object in array
end


////////////////////
////////////////////
//*) make a class w/ random variable
//*) randomize it
//*) now, randomize just one of the members of the class.
//*) add a constraint. Do the same




   


