// Stand-alone test inside program block
program testcase(//Inputs to Design, Outputs from Program <-- Signals are to be driven inside Progam Block

                 //Inout to/from Design, inout to/from Programa <-- Signals are to be driven inside Program

                 //Output from Design, Input to Program <-- Signals are to be monitored

                );

   initial begin
      ...
   end

endprogram
