module testbench();



endmodule
