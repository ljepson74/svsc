class packet;
   
   // your code here
endclass
