module top;
   initial begin

      $display("start---------");

      $display("one two \
3three");
   end


endmodule
