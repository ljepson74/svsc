module top;


endmodule