library ieee;   
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity my_vhdl is
  port (
    bus : in std_logic_vector(3 downto 0);
  );

end my_vhdl;

--architecture arch of my_vhdl is
--
--begin  -- arch
--
--  
--
--end arch;
