module q();

   initial begin
      repeat (5) $display("************** THIS WORKED. *******");
   end
   
endmodule