// TITLE: Some other title

// Presence of this comment here causes the below class to get missed.
// Class: MISS1
// this will get missed, I think, b/c line above Class:

// CLASS: TOP2
// This is my second class code.  CLASS and Class both work btw.  IMG MIPS is pushing we uniformly use "CLASS"

 class top2();

// VARIABLE: fred
   int fred;
      
// VARIABLE: red

   int red;

// VARIABLE:
   int red1;
   int red2;
   int red3;

      
endclass

// Class: MISS2
// this will not get missed, I think
