interface c_if(
		   input clk
		   );
   logic 		 my_signal;

endinterface // c_if

