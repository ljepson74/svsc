class kl_class;
    function void whoami(input string name="hossein");
       $display("my name is %0s",name);
    endfunction : whoami
endclass // kl_class
