//this is a basic class

class class_abc; 
   rand int n1;
   rand int n2;     
endclass // abc

