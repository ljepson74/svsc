
task init();
  reset = 1;
  enable = 0;
  preload = 0;
  mode = 0;
endtask
