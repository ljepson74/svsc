class c1;
   c2 my_c2;
   
   
   function new();      
      $display(" %m: MADE C1");      
      my_c2  = new();      
   endfunction // new
   
endclass // c1
