package iclp_pkg;
  //plusargs are bit(a boolean), an int, or a string
   typedef enum {BIT=0, INT=1, STRING=2} valuetype_e;  //this is now defined twice
endpackage : iclp_pkg
   