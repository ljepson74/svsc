

module top();


   mod_wants_assoc_array  mod_wants_assoc_array();
   mod_w_assoc_array      mod_w_assoc_array();

endmodule // top

  
