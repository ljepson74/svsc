module top_level;

   access_other_modules_data_play access_other_modules_data_play();

   other_module other_module();

endmodule // top_level
