// PACKAGE: package1

package package1;

endpackage // package1
   