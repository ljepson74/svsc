// FRIENDSHIP: horse
class horse();
endclass // horse
